.title KiCad schematic
R11 +5V Net-_NMOS16-D_ R_Small
NMOS16 __NMOS16
R0 +5V Net-_NMOS0-D_ R_Small
NMOS0 __NMOS0
NMOS6 __NMOS6
R5 +5V Net-_NMOS15-G_ R_Small
R2 +5V Net-_NMOS2-D_ R_Small
NMOS2 __NMOS2
NMOS3 __NMOS3
NMOS1 __NMOS1
R1 +5V Net-_NMOS1-D_ R_Small
R9 +5V Net-_NMOS14-D_ R_Small
NMOS14 __NMOS14
R10 +5V Net-_NMOS15-D_ R_Small
NMOS15 __NMOS15
R13 +5V /CTRL4 R_Small
NMOS18 __NMOS18
NMOS19 __NMOS19
R12 +5V Net-_NMOS17-D_ R_Small
NMOS17 __NMOS17
NMOS7 __NMOS7
NMOS8 __NMOS8
R6 +5V /CTRL5 R_Small
NMOS9 __NMOS9
NMOS10 __NMOS10
R7 +5V Net-_NMOS10-D_ R_Small
NMOS11 __NMOS11
R4 +5V Net-_NMOS10-G_ R_Small
NMOS5 __NMOS5
R3 +5V Net-_NMOS11-G_ R_Small
NMOS4 __NMOS4
R8 +5V /CTRL8 R_Small
NMOS12 __NMOS12
NMOS13 __NMOS13
.end
